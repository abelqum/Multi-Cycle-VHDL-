library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity RAM is
port(
    clk     : in  std_logic; 
    Adress  : in  std_logic_vector(7 downto 0);
    Data_in : in  std_logic_vector(23 downto 0);
    EnRAM   : in  std_logic; 
    RW      : in  std_logic; 
    Data_out: out std_logic_vector(23 downto 0)
);
end RAM;

architecture Behavioral of RAM is

   type RAM_MEMORY is array (0 to 255) of std_logic_vector(23 downto 0);

signal MEMORY: RAM_MEMORY := (
    -- PROGRAMA 1: 17x+25y-w/4
    -- W=27 (en 217), X=3 (en 218), Y=15 (en 219)
    0 => "00001011" & "00000000" & "11011000",  -- LW R0, [W] (Offset=216 -> PC+1+Off = 1+216=217)
    1 => "00001011" & "00000001" & "11011000",  -- LW R1, [X] (Offset=216 -> PC+1+Off = 2+216=218)
    2 => "00001011" & "00000010" & "11011000",  -- LW R2, [Y] (Offset=216 -> PC+1+Off = 3+216=219)
    
    -- Calcular 17X
    3 => "00011101" & "00000001" & "00010001",  -- MULI R1, 17 (R1 = 3 * 17 = 51)
    4 => "00100101" & "00000001" & "00000000",  -- DISP R1 (Muestra 51)
    
    -- Calcular 25Y    
    5 => "00011101" & "00000010" & "00011001",  -- MULI R2, 25 (R2 = 15 * 25 = 375)
    6 => "00100101" & "00000010" & "00000000",  -- DISP R2 (Muestra 375)
    
    -- Calcular W/4
    7 => "00011110" & "00000000" & "00000100",  -- DIVI R0, 4 (R0 = 27 / 4 = 6)
    8 => "00100101" & "00000000" & "00000000",  -- DISP R0 (Muestra 6)
    
    -- Calcular 17X + 25Y
    9 => "00000000" & "00000001" & "00000010",  -- ADD R1, R2 (R1 = 51 + 375 = 426)
    10 => "00100101" & "00000001" & "00000000", -- DISP R1 (Muestra 426)
    
    -- Calcular (17X + 25Y) - W/4 
    11 => "00000001" & "00000001" & "00000000", -- SUB R1, R0 (R1 = 426 - 6 = 420)
    12 => "00100101" & "00000001" & "00000000", -- DISP R1 (Muestra 420)
    
    13 => "00100100" & "00000000" & "00000000", -- HALT 

    -- FIN PROGRAMA 1

    
    -- PROGRAMA 2: 10x^2 + 30x - z/2
    -- Inicia en 14. X=3 (en 218), Z=19 (en 220)
    14 => "00001011" & "00000000" & "11001011", -- LW R0, [X] (Offset=203 -> PC+1+Off = 15+203=218)
    15 => "00001011" & "00000001" & "11001010", -- LW R1, [X] (Offset=202 -> PC+1+Off = 16+202=218)
    16 => "00001011" & "00000010" & "11001100", -- LW R2, [Z] (Offset=204 -> PC+1+Off = 17+204=220)
    
    -- Calcular X^2 (X * X)
    17 => "00000010" & "00000000" & "00000000", -- MUL R0, R0  (R0 = 3 * 3 = 9)
    18 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 9)
    
    -- Calcular 10X^2 (Sobrescribe R0)
    19 => "00011101" & "00000000" & "00001010", -- MULI R0, 10 (R0 = 9 * 10 = 90)
    20 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 90)
    
    -- Calcular 30X
    21 => "00011101" & "00000001" & "00011110", -- MULI R1, 30 (R1 = 3 * 30 = 90) 
    22 => "00100101" & "00000001" & "00000000", -- DISP R1 (Muestra 90)
    
    -- Sumar 10X^2 + 30X
    23 => "00000000" & "00000000" & "00000001", -- ADD R0, R1 (R0 = 90 + 90 = 180)
    24 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 180)
    
    -- Calcular Z/2
    25 => "00011110" & "00000010" & "00000010", -- DIVI R2, 2 (R2 = 19 / 2 = 9)
    26 => "00100101" & "00000010" & "00000000", -- DISP R2 (Muestra 9)
    
    -- Calcular (10X^2 + 30X) - Z/2
    27 => "00000001" & "00000000" & "00000010", -- SUB R0, R2 (R0 = 180 - 9 = 171)
    28 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 171)
    
    29 => "00100100" & "00000000" & "00000000", -- HALT 
      -- FIN PROGRAMA 2


    -- PROGRAMA 3: -X^3 – 7Z+ W / (10)
    -- Inicia en 30. W=27 (en 217), X=3 (en 218), Z=19 (en 220)
    30 => "00001011" & "00000000" & "10111010", -- LW R0, [W] (Offset=186 -> PC+1+Off = 31+186=217)
    31 => "00001011" & "00000001" & "10111010", -- LW R1, [X] (Offset=186 -> PC+1+Off = 32+186=218)
    32 => "00001011" & "00000010" & "10111011", -- LW R2, [Z] (Offset=187 -> PC+1+Off = 33+187=220)
    33 => "00001011" & "00000011" & "10111000", -- LW R3, [X] (Offset=184 -> PC+1+Off = 34+184=218)
    
    34 => "00000010" & "00000001" & "00000001", -- MUL R1, R1 (R1 = 3 * 3 = 9) (X^2)
    35 => "00100101" & "00000001" & "00000000", -- DISP R1 (Muestra 9)
    
    36 => "00000010" & "00000001" & "00000011", -- MUL R1, R3 (R1 = 9 * 3 = 27) (X^3)
    37 => "00100101" & "00000001" & "00000000", -- DISP R1 (Muestra 27)
    
    38 => "00011101" & "00000010" & "00000111", -- MULI R2, 7 (R2 = 19 * 7 = 133) (7Z)
    39 => "00100101" & "00000010" & "00000000", -- DISP R2 (Muestra 133)
    
    40 => "00011110" & "00000000" & "00001010", -- DIVI R0, 10 (R0 = 27 / 10 = 2) (W/10)
    41 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 2)
    
    42 => "00000001" & "00000000" & "00000010", -- SUB R0, R2 (R0 = 2 - 133 = -131)
    43 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra -131)
    
    44 => "00000001" & "00000000" & "00000001", -- SUB R0, R1 (R0 = -131 - 27 = -158)
    45 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra -158)
    
    46 => "00100100" & "00000000" & "00000000", -- HALT 
    -- FIN PROGRAMA 3

    -- PROGRAMA 4
    47 => "00100100" & "00000000" & "00000000",  -- HALT
    -- FIN PROGRAMA 4

    -- =================================================================
    -- PROGRAMA 5 (PRACTICA 2A - SIN DELAYS)
    -- Inicia en 48. DATOS en 221-230
    -- =================================================================
    -- R0=Dato, R2=Zero, R3=Imm
    48 => "00000001" & "00000010" & "00000010", -- SUB R2, R2 (R2 = 0, 'Zero')

    -- === Bloque 1: W (1003) @221 + 5 ===
    49 => "00001011" & "00000000" & "10101011", -- LW R0, [W_P2A] (Offset=171 -> PC+1+Off = 50+171=221)
    50 => "00011011" & "00000011" & "00000101", -- ADDI R3, R2, 5 (R3 = 5)
    51 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 1003 + 5 = 1008)
    52 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 1008)

    -- === Bloque 2: X (101) @222 + 6 ===
    53 => "00001011" & "00000000" & "10101000", -- LW R0, [X_P2A] (Offset=168 -> PC+1+Off = 54+168=222)
    54 => "00011011" & "00000011" & "00000110", -- ADDI R3, R2, 6 (R3 = 6)
    55 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 101 + 6 = 107)
    56 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 107)

    -- === Bloque 3: Y (70) @223 + 7 ===
    57 => "00001011" & "00000000" & "10100101", -- LW R0, [Y_P2A] (Offset=165 -> PC+1+Off = 58+165=223)
    58 => "00011011" & "00000011" & "00000111", -- ADDI R3, R2, 7 (R3 = 7)
    59 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 70 + 7 = 77)
    60 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 77)

    -- === Bloque 4: Z (50) @224 + 8 ===
    61 => "00001011" & "00000000" & "10100010", -- LW R0, [Z_P2A] (Offset=162 -> PC+1+Off = 62+162=224)
    62 => "00011011" & "00000011" & "00001000", -- ADDI R3, R2, 8 (R3 = 8)
    63 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 50 + 8 = 58)
    64 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 58)

    -- === Bloque 5: M (18) @225 + 9 ===
    65 => "00001011" & "00000000" & "10011111", -- LW R0, [M_P2A] (Offset=159 -> PC+1+Off = 66+159=225)
    66 => "00011011" & "00000011" & "00001001", -- ADDI R3, R2, 9 (R3 = 9)
    67 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 18 + 9 = 27)
    68 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 27)

    -- === Bloque 6: N (7) @226 + 10 ===
    69 => "00001011" & "00000000" & "10011100", -- LW R0, [N_P2A] (Offset=156 -> PC+1+Off = 70+156=226)
    70 => "00011011" & "00000011" & "00001010", -- ADDI R3, R2, 10 (R3 = 10)
    71 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 7 + 10 = 17)
    72 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 17)
    
    -- === Bloque 7: O (23) @227 + 11 ===
    73 => "00001011" & "00000000" & "10011001", -- LW R0, [O_P2A] (Offset=153 -> PC+1+Off = 74+153=227)
    74 => "00011011" & "00000011" & "00001011", -- ADDI R3, R2, 11 (R3 = 11)
    75 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 23 + 11 = 34)
    76 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 34)

    -- === Bloque 8: P (55) @228 + 12 ===
    77 => "00001011" & "00000000" & "10010110", -- LW R0, [P_P2A] (Offset=150 -> PC+1+Off = 78+150=228)
    78 => "00011011" & "00000011" & "00001100", -- ADDI R3, R2, 12 (R3 = 12)
    79 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 55 + 12 = 67)
    80 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 67)

    -- === Bloque 9: Q (77) @229 + 13 ===
    81 => "00001011" & "00000000" & "10010011", -- LW R0, [Q_P2A] (Offset=147 -> PC+1+Off = 82+147=229)
    82 => "00011011" & "00000011" & "00001101", -- ADDI R3, R2, 13 (R3 = 13)
    83 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 77 + 13 = 90)
    84 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 90)

    -- === Bloque 10: R (19) @230 + 14 ===
    85 => "00001011" & "00000000" & "10010000", -- LW R0, [R_P2A] (Offset=144 -> PC+1+Off = 86+144=230)
    86 => "00011011" & "00000011" & "00001110", -- ADDI R3, R2, 14 (R3 = 14)
    87 => "00000000" & "00000000" & "00000011", -- ADD R0, R3 (R0 = 19 + 14 = 33)
    88 => "00100101" & "00000000" & "00000000", -- DISP R0 (Muestra 33)

    -- FIN PROGRAMA 5
    89 => "00100100" & "00000000" & "00000000", -- HALT


    -- ... (Espacio vacío)


    -- =================================================================
    -- SECCIÓN DE DATOS (A partir de 217, como en tu código)
    -- =================================================================
    217 => "00000000" & "00000000" & "00011011",  -- W = 27 decimal
    218 => "00000000" & "00000000" & "00000011",  -- X = 3 decimal
    219 => "00000000" & "00000000" & "00001111",  -- Y = 15 decimal
    220 => "00000000" & "00000000" & "00010011",  -- Z = 19 decimal
    --SECCIÓN DE DATOS PRÁCTICA 2
    221 => "00000000" & "00000011" & "11101011",  -- W_P2A = 1003
    222 => "00000000" & "00000000" & "01100101",  -- X_P2A = 101
    223 => "00000000" & "00000000" & "01000110",  -- Y_P2A = 70
    224 => "00000000" & "00000000" & "00110010",  -- Z_P2A = 50
    225 => "00000000" & "00000000" & "00010010",  -- M_P2A = 18
    226 => "00000000" & "00000000" & "00000111",  -- N_P2A = 7
    227 => "00000000" & "00000000" & "00010111",  -- O_P2A = 23
    228 => "00000000" & "00000000" & "00110111",  -- P_P2A = 55
    229 => "00000000" & "00000000" & "01001101",  -- Q_P2A = 77
    230 => "00000000" & "00000000" & "00010011",  -- R_P2A = 19
    
    others => (others => '0')
);
  signal addr_int : integer range 0 to 255; 
--    
begin
 
    addr_int <= to_integer(unsigned(Adress));

    -- Escritura Síncrona
    process(clk)
    begin
        if rising_edge(clk) then
            if EnRAM = '1' and RW = '0' then 
                MEMORY(addr_int) <= Data_in; 
            end if;
        end if;
    end process;

    -- Lectura Asíncrona
    Data_out <= MEMORY(addr_int);

end Behavioral;
