library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity RAM is
port(
    clk     : in  std_logic; 
    Adress  : in  std_logic_vector(7 downto 0);
    Data_in : in  std_logic_vector(23 downto 0);
    EnRAM   : in  std_logic; 
    RW      : in  std_logic; 
    Data_out: out std_logic_vector(23 downto 0)
);
end RAM;

architecture Behavioral of RAM is

   type RAM_MEMORY is array (0 to 255) of std_logic_vector(23 downto 0);

signal RAM_array : RAM_type := (
    -- ============ ECUACIÓN A: F(X,Y,W) = 17X + 25Y - W/4 ============
    -- Asumiendo: X en RF@1, Y en RF@2, W en RF@3
    0   => "00001011" & "00000001" & "00000000",  -- MOVRR RF@1 -> RF@0 (X)
    1   => "00011100" & "00000000" & "00010000",  -- LSLI RF@0, 4 (X*16)  
    2   => "00011011" & "00000001" & "00010000",  -- MOVRR RF@1 -> RF@4 (copia X)
    3   => "00000000" & "00000000" & "00010000",  -- ADD RF@0, RF@4 (16X+X=17X)
    4   => "00011011" & "00000010" & "00010101",  -- MOVRR RF@2 -> RF@5 (Y)
    5   => "00011100" & "00000101" & "00010000",  -- LSLI RF@5, 4 (Y*16)
    6   => "00011011" & "00000010" & "00010110",  -- MOVRR RF@2 -> RF@6 (copia Y)
    7   => "00011100" & "00000110" & "00011000",  -- LSLI RF@6, 3 (Y*8)
    8   => "00000000" & "00000101" & "00010110",  -- ADD RF@5, RF@6 (16Y+8Y)
    9   => "00011011" & "00000010" & "00010111",  -- MOVRR RF@2 -> RF@7 (copia Y)
    10  => "00000000" & "00000101" & "00010111",  -- ADD RF@5, RF@7 (+Y = 25Y)
    11  => "00000000" & "00000000" & "00010101",  -- ADD RF@0, RF@5 (17X+25Y)
    12  => "00011011" & "00000011" & "00010110",  -- MOVRR RF@3 -> RF@6 (W)
    13  => "00011101" & "00000110" & "00000010",  -- ASRI RF@6, 2 (W/4)
    14  => "00000001" & "00000000" & "00010110",  -- SUB RF@0, RF@6 (result-W/4)
    15  => "00100100" & "00000000" & "00000000",  -- HALT

    -- ============ ECUACIÓN B: F(X,Z) = 10X² + 30X - Z/2 ============
    -- Asumiendo: X en RF@1, Z en RF@4
    32  => "00011011" & "00000001" & "00000000",  -- MOVRR RF@1 -> RF@0 (X)
    33  => "00000010" & "00000000" & "00000000",  -- MULT RF@0, RF@0 (X²)
    34  => "00011011" & "00000000" & "00010001",  -- MOVRR RF@0 -> RF@1 (copia X²)
    35  => "00011100" & "00000001" & "00011000",  -- LSLI RF@1, 3 (8X²)
    36  => "00011011" & "00000000" & "00010010",  -- MOVRR RF@0 -> RF@2 (copia X²)
    37  => "00011100" & "00000010" & "00010000",  -- LSLI RF@2, 1 (2X²)
    38  => "00000000" & "00000001" & "00010010",  -- ADD RF@1, RF@2 (10X²)
    39  => "00011011" & "00000001" & "00010011",  -- MOVRR RF@1 -> RF@3 (copia X)
    40  => "00011100" & "00000011" & "00100000",  -- LSLI RF@3, 4 (16X)
    41  => "00011011" & "00000001" & "00010100",  -- MOVRR RF@1 -> RF@4 (copia X)
    42  => "00011100" & "00000100" & "00011000",  -- LSLI RF@4, 3 (8X)
    43  => "00000000" & "00000011" & "00010100",  -- ADD RF@3, RF@4 (16X+8X)
    44  => "00011011" & "00000001" & "00010101",  -- MOVRR RF@1 -> RF@5 (copia X)
    45  => "00011100" & "00000101" & "00010000",  -- LSLI RF@5, 2 (4X)
    46  => "00000000" & "00000011" & "00010101",  -- ADD RF@3, RF@5 (+4X)
    47  => "00011011" & "00000001" & "00010110",  -- MOVRR RF@1 -> RF@6 (copia X)
    48  => "00011100" & "00000110" & "00010000",  -- LSLI RF@6, 1 (2X)
    49  => "00000000" & "00000011" & "00010110",  -- ADD RF@3, RF@6 (+2X = 30X)
    50  => "00000000" & "00000001" & "00010011",  -- ADD RF@1, RF@3 (10X²+30X)
    51  => "00011011" & "00000100" & "00010111",  -- MOVRR RF@4 -> RF@7 (Z)
    52  => "00011101" & "00000111" & "00000001",  -- ASRI RF@7, 1 (Z/2)
    53  => "00000001" & "00000001" & "00010111",  -- SUB RF@1, RF@7 (result-Z/2)
    54  => "00100100" & "00000000" & "00000000",  -- HALT

    -- ============ ECUACIÓN C: F(X,Z,W) = -X³ - 7Z + W/10 ============
    -- Asumiendo: X en RF@1, Z en RF@4, W en RF@5
    64  => "00011011" & "00000001" & "00000000",  -- MOVRR RF@1 -> RF@0 (X)
    65  => "00000010" & "00000000" & "00000000",  -- MULT RF@0, RF@0 (X²)
    66  => "00000010" & "00000000" & "00000001",  -- MULT RF@0, RF@1 (X³)
    67  => "00000111" & "00000000" & "00000000",  -- COMP1 RF@0 (comp1 X³)
    68  => "00001000" & "00000000" & "00000000",  -- COMP2 RF@0 (-X³)
    69  => "00011011" & "00000100" & "00010001",  -- MOVRR RF@4 -> RF@1 (Z)
    70  => "00011100" & "00000001" & "00010000",  -- LSLI RF@1, 2 (4Z)
    71  => "00011011" & "00000100" & "00010010",  -- MOVRR RF@4 -> RF@2 (copia Z)
    72  => "00011100" & "00000010" & "00010000",  -- LSLI RF@2, 1 (2Z)
    73  => "00000000" & "00000001" & "00010010",  -- ADD RF@1, RF@2 (4Z+2Z)
    74  => "00011011" & "00000100" & "00010011",  -- MOVRR RF@4 -> RF@3 (copia Z)
    75  => "00000000" & "00000001" & "00010011",  -- ADD RF@1, RF@3 (+Z = 7Z)
    76  => "00000001" & "00000000" & "00010001",  -- SUB RF@0, RF@1 (-X³-7Z)
    77  => "00011011" & "00000101" & "00010100",  -- MOVRR RF@5 -> RF@4 (W)
    78  => "00011101" & "00000100" & "00000011",  -- ASRI RF@4, 3 (W/8)
    79  => "00011011" & "00000101" & "00010101",  -- MOVRR RF@5 -> RF@5 (copia W)
    80  => "00011101" & "00000101" & "00000101",  -- ASRI RF@5, 5 (W/32)
    81  => "00000000" & "00000100" & "00010101",  -- ADD RF@4, RF@5 (W/8+W/32≈W/10)
    82  => "00000000" & "00000000" & "00010100",  -- ADD RF@0, RF@4 (result+W/10)
    83  => "00100100" & "00000000" & "00000000",  -- HALT

    -- ============ ECUACIÓN D: Desplegar "0000" ============
    96  => "00011011" & "00000000" & "00000000",  -- MOVRR RF@0 -> RF@0 (0)
    97  => "00011011" & "00000000" & "00010001",  -- MOVRR RF@0 -> RF@1 (0)
    98  => "00011011" & "00000000" & "00010010",  -- MOVRR RF@0 -> RF@2 (0)
    99  => "00011011" & "00000000" & "00010011",  -- MOVRR RF@0 -> RF@3 (0)
    100 => "00011011" & "00000000" & "00010100",  -- MOVRR RF@0 -> RF@4 (0)
    101 => "00100100" & "00000000" & "00000000",  -- HALT

    others => "00000000" & "00000000" & "00000000"
);
  signal addr_int : integer range 0 to 255; 

begin

    addr_int <= to_integer(unsigned(Adress));

    -- Escritura Síncrona
    process(clk)
    begin
        if rising_edge(clk) then
            if EnRAM = '1' and RW = '0' then 
                MEMORY(addr_int) <= Data_in; 
            end if;
        end if;
    end process;

    -- Lectura Asíncrona
    Data_out <= MEMORY(addr_int);

end Behavioral;